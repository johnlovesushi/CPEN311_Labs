-- DE1_SoC_QSYS_audio.vhd

-- Generated using ACDS version 14.1 186 at 2017.11.28.14:38:56

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE1_SoC_QSYS_audio is
	port (
		clk_clk                      : in  std_logic                     := '0';             --               clk.clk
		data_divfrec_export          : out std_logic_vector(31 downto 0);                    --      data_divfrec.export
		data_fregen_s1_address       : in  std_logic_vector(1 downto 0)  := (others => '0'); --    data_fregen_s1.address
		data_fregen_s1_write_n       : in  std_logic                     := '0';             --                  .write_n
		data_fregen_s1_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		data_fregen_s1_chipselect    : in  std_logic                     := '0';             --                  .chipselect
		data_fregen_s1_readdata      : out std_logic_vector(31 downto 0);                    --                  .readdata
		empty_export                 : in  std_logic                     := '0';             --             empty.export
		empty_s1_address             : in  std_logic_vector(1 downto 0)  := (others => '0'); --          empty_s1.address
		empty_s1_readdata            : out std_logic_vector(31 downto 0);                    --                  .readdata
		fifo_full_export             : in  std_logic                     := '0';             --         fifo_full.export
		fifo_full_s1_address         : in  std_logic_vector(1 downto 0)  := (others => '0'); --      fifo_full_s1.address
		fifo_full_s1_readdata        : out std_logic_vector(31 downto 0);                    --                  .readdata
		fifo_used_export             : in  std_logic_vector(11 downto 0) := (others => '0'); --         fifo_used.export
		fifo_used_s1_address         : in  std_logic_vector(1 downto 0)  := (others => '0'); --      fifo_used_s1.address
		fifo_used_s1_readdata        : out std_logic_vector(31 downto 0);                    --                  .readdata
		out_data_audio_export        : out std_logic_vector(31 downto 0);                    --    out_data_audio.export
		out_data_audio_s1_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- out_data_audio_s1.address
		out_data_audio_s1_write_n    : in  std_logic                     := '0';             --                  .write_n
		out_data_audio_s1_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		out_data_audio_s1_chipselect : in  std_logic                     := '0';             --                  .chipselect
		out_data_audio_s1_readdata   : out std_logic_vector(31 downto 0);                    --                  .readdata
		out_pause_export             : out std_logic;                                        --         out_pause.export
		out_pause_s1_address         : in  std_logic_vector(1 downto 0)  := (others => '0'); --      out_pause_s1.address
		out_pause_s1_write_n         : in  std_logic                     := '0';             --                  .write_n
		out_pause_s1_writedata       : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		out_pause_s1_chipselect      : in  std_logic                     := '0';             --                  .chipselect
		out_pause_s1_readdata        : out std_logic_vector(31 downto 0);                    --                  .readdata
		out_stop_export              : out std_logic;                                        --          out_stop.export
		out_stop_s1_address          : in  std_logic_vector(1 downto 0)  := (others => '0'); --       out_stop_s1.address
		out_stop_s1_write_n          : in  std_logic                     := '0';             --                  .write_n
		out_stop_s1_writedata        : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		out_stop_s1_chipselect       : in  std_logic                     := '0';             --                  .chipselect
		out_stop_s1_readdata         : out std_logic_vector(31 downto 0);                    --                  .readdata
		reset_reset_n                : in  std_logic                     := '0';             --             reset.reset_n
		wrclk_export                 : out std_logic;                                        --             wrclk.export
		wrclk_s1_address             : in  std_logic_vector(1 downto 0)  := (others => '0'); --          wrclk_s1.address
		wrclk_s1_write_n             : in  std_logic                     := '0';             --                  .write_n
		wrclk_s1_writedata           : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		wrclk_s1_chipselect          : in  std_logic                     := '0';             --                  .chipselect
		wrclk_s1_readdata            : out std_logic_vector(31 downto 0);                    --                  .readdata
		wrreq_export                 : out std_logic;                                        --             wrreq.export
		wrreq_s1_address             : in  std_logic_vector(1 downto 0)  := (others => '0'); --          wrreq_s1.address
		wrreq_s1_write_n             : in  std_logic                     := '0';             --                  .write_n
		wrreq_s1_writedata           : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		wrreq_s1_chipselect          : in  std_logic                     := '0';             --                  .chipselect
		wrreq_s1_readdata            : out std_logic_vector(31 downto 0)                     --                  .readdata
	);
end entity DE1_SoC_QSYS_audio;

architecture rtl of DE1_SoC_QSYS_audio is
	component DE1_SoC_QSYS_audio_DATA_FREGEN is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component DE1_SoC_QSYS_audio_DATA_FREGEN;

	component DE1_SoC_QSYS_audio_EMPTY is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component DE1_SoC_QSYS_audio_EMPTY;

	component DE1_SoC_QSYS_audio_OUT_PAUSE is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component DE1_SoC_QSYS_audio_OUT_PAUSE;

	component DE1_SoC_QSYS_audio_fifo_used is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(11 downto 0) := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_audio_fifo_used;

begin

	data_fregen : component DE1_SoC_QSYS_audio_DATA_FREGEN
		port map (
			clk        => clk_clk,                   --                 clk.clk
			reset_n    => reset_reset_n,             --               reset.reset_n
			address    => data_fregen_s1_address,    --                  s1.address
			write_n    => data_fregen_s1_write_n,    --                    .write_n
			writedata  => data_fregen_s1_writedata,  --                    .writedata
			chipselect => data_fregen_s1_chipselect, --                    .chipselect
			readdata   => data_fregen_s1_readdata,   --                    .readdata
			out_port   => data_divfrec_export        -- external_connection.export
		);

	empty : component DE1_SoC_QSYS_audio_EMPTY
		port map (
			clk      => clk_clk,           --                 clk.clk
			reset_n  => reset_reset_n,     --               reset.reset_n
			address  => empty_s1_address,  --                  s1.address
			readdata => empty_s1_readdata, --                    .readdata
			in_port  => empty_export       -- external_connection.export
		);

	fifo_full : component DE1_SoC_QSYS_audio_EMPTY
		port map (
			clk      => clk_clk,               --                 clk.clk
			reset_n  => reset_reset_n,         --               reset.reset_n
			address  => fifo_full_s1_address,  --                  s1.address
			readdata => fifo_full_s1_readdata, --                    .readdata
			in_port  => fifo_full_export       -- external_connection.export
		);

	out_data_audio : component DE1_SoC_QSYS_audio_DATA_FREGEN
		port map (
			clk        => clk_clk,                      --                 clk.clk
			reset_n    => reset_reset_n,                --               reset.reset_n
			address    => out_data_audio_s1_address,    --                  s1.address
			write_n    => out_data_audio_s1_write_n,    --                    .write_n
			writedata  => out_data_audio_s1_writedata,  --                    .writedata
			chipselect => out_data_audio_s1_chipselect, --                    .chipselect
			readdata   => out_data_audio_s1_readdata,   --                    .readdata
			out_port   => out_data_audio_export         -- external_connection.export
		);

	out_pause : component DE1_SoC_QSYS_audio_OUT_PAUSE
		port map (
			clk        => clk_clk,                 --                 clk.clk
			reset_n    => reset_reset_n,           --               reset.reset_n
			address    => out_pause_s1_address,    --                  s1.address
			write_n    => out_pause_s1_write_n,    --                    .write_n
			writedata  => out_pause_s1_writedata,  --                    .writedata
			chipselect => out_pause_s1_chipselect, --                    .chipselect
			readdata   => out_pause_s1_readdata,   --                    .readdata
			out_port   => out_pause_export         -- external_connection.export
		);

	out_stop : component DE1_SoC_QSYS_audio_OUT_PAUSE
		port map (
			clk        => clk_clk,                --                 clk.clk
			reset_n    => reset_reset_n,          --               reset.reset_n
			address    => out_stop_s1_address,    --                  s1.address
			write_n    => out_stop_s1_write_n,    --                    .write_n
			writedata  => out_stop_s1_writedata,  --                    .writedata
			chipselect => out_stop_s1_chipselect, --                    .chipselect
			readdata   => out_stop_s1_readdata,   --                    .readdata
			out_port   => out_stop_export         -- external_connection.export
		);

	wrclk : component DE1_SoC_QSYS_audio_OUT_PAUSE
		port map (
			clk        => clk_clk,             --                 clk.clk
			reset_n    => reset_reset_n,       --               reset.reset_n
			address    => wrclk_s1_address,    --                  s1.address
			write_n    => wrclk_s1_write_n,    --                    .write_n
			writedata  => wrclk_s1_writedata,  --                    .writedata
			chipselect => wrclk_s1_chipselect, --                    .chipselect
			readdata   => wrclk_s1_readdata,   --                    .readdata
			out_port   => wrclk_export         -- external_connection.export
		);

	wrreq : component DE1_SoC_QSYS_audio_OUT_PAUSE
		port map (
			clk        => clk_clk,             --                 clk.clk
			reset_n    => reset_reset_n,       --               reset.reset_n
			address    => wrreq_s1_address,    --                  s1.address
			write_n    => wrreq_s1_write_n,    --                    .write_n
			writedata  => wrreq_s1_writedata,  --                    .writedata
			chipselect => wrreq_s1_chipselect, --                    .chipselect
			readdata   => wrreq_s1_readdata,   --                    .readdata
			out_port   => wrreq_export         -- external_connection.export
		);

	fifo_used : component DE1_SoC_QSYS_audio_fifo_used
		port map (
			clk      => clk_clk,               --                 clk.clk
			reset_n  => reset_reset_n,         --               reset.reset_n
			address  => fifo_used_s1_address,  --                  s1.address
			readdata => fifo_used_s1_readdata, --                    .readdata
			in_port  => fifo_used_export       -- external_connection.export
		);

end architecture rtl; -- of DE1_SoC_QSYS_audio
