-- DE1_SoC_QSYS.vhd

-- Generated using ACDS version 14.1 186 at 2017.11.28.14:38:55

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE1_SoC_QSYS is
	port (
		audio2fifo_0_data_divfrec_export                  : out   std_logic_vector(31 downto 0);                    --                  audio2fifo_0_data_divfrec.export
		audio2fifo_0_empty_export                         : in    std_logic                     := '0';             --                         audio2fifo_0_empty.export
		audio2fifo_0_fifo_full_export                     : in    std_logic                     := '0';             --                     audio2fifo_0_fifo_full.export
		audio2fifo_0_fifo_used_export                     : in    std_logic_vector(11 downto 0) := (others => '0'); --                     audio2fifo_0_fifo_used.export
		audio2fifo_0_out_data_audio_export                : out   std_logic_vector(31 downto 0);                    --                audio2fifo_0_out_data_audio.export
		audio2fifo_0_out_pause_export                     : out   std_logic;                                        --                     audio2fifo_0_out_pause.export
		audio2fifo_0_out_stop_export                      : out   std_logic;                                        --                      audio2fifo_0_out_stop.export
		audio2fifo_0_wrclk_export                         : out   std_logic;                                        --                         audio2fifo_0_wrclk.export
		audio2fifo_0_wrreq_export                         : out   std_logic;                                        --                         audio2fifo_0_wrreq.export
		audio_sel_export                                  : out   std_logic;                                        --                                  audio_sel.export
		clk_clk                                           : in    std_logic                     := '0';             --                                        clk.clk
		clk_25_out_clk                                    : out   std_logic;                                        --                                 clk_25_out.clk
		clk_sdram_clk                                     : out   std_logic;                                        --                                  clk_sdram.clk
		dds_increment_external_connection_export          : out   std_logic_vector(31 downto 0);                    --          dds_increment_external_connection.export
		div_freq_export                                   : out   std_logic_vector(31 downto 0);                    --                                   div_freq.export
		key_external_connection_export                    : in    std_logic_vector(3 downto 0)  := (others => '0'); --                    key_external_connection.export
		keyboard_keys_export                              : in    std_logic_vector(31 downto 0) := (others => '0'); --                              keyboard_keys.export
		lfsr_clk_interrupt_gen_external_connection_export : in    std_logic                     := '0';             -- lfsr_clk_interrupt_gen_external_connection.export
		lfsr_val_external_connection_export               : in    std_logic_vector(31 downto 0) := (others => '0'); --               lfsr_val_external_connection.export
		modulation_selector_export                        : out   std_logic_vector(3 downto 0);                     --                        modulation_selector.export
		mouse_pos_export                                  : in    std_logic_vector(31 downto 0) := (others => '0'); --                                  mouse_pos.export
		pll_locked_export                                 : out   std_logic;                                        --                                 pll_locked.export
		reset_reset_n                                     : in    std_logic                     := '0';             --                                      reset.reset_n
		sdram_wire_addr                                   : out   std_logic_vector(12 downto 0);                    --                                 sdram_wire.addr
		sdram_wire_ba                                     : out   std_logic_vector(1 downto 0);                     --                                           .ba
		sdram_wire_cas_n                                  : out   std_logic;                                        --                                           .cas_n
		sdram_wire_cke                                    : out   std_logic;                                        --                                           .cke
		sdram_wire_cs_n                                   : out   std_logic;                                        --                                           .cs_n
		sdram_wire_dq                                     : inout std_logic_vector(15 downto 0) := (others => '0'); --                                           .dq
		sdram_wire_dqm                                    : out   std_logic_vector(1 downto 0);                     --                                           .dqm
		sdram_wire_ras_n                                  : out   std_logic;                                        --                                           .ras_n
		sdram_wire_we_n                                   : out   std_logic;                                        --                                           .we_n
		signal_selector_export                            : out   std_logic_vector(7 downto 0);                     --                            signal_selector.export
		vga_alt_vip_itc_0_clocked_video_vid_clk           : in    std_logic                     := '0';             --            vga_alt_vip_itc_0_clocked_video.vid_clk
		vga_alt_vip_itc_0_clocked_video_vid_data          : out   std_logic_vector(23 downto 0);                    --                                           .vid_data
		vga_alt_vip_itc_0_clocked_video_underflow         : out   std_logic;                                        --                                           .underflow
		vga_alt_vip_itc_0_clocked_video_vid_datavalid     : out   std_logic;                                        --                                           .vid_datavalid
		vga_alt_vip_itc_0_clocked_video_vid_v_sync        : out   std_logic;                                        --                                           .vid_v_sync
		vga_alt_vip_itc_0_clocked_video_vid_h_sync        : out   std_logic;                                        --                                           .vid_h_sync
		vga_alt_vip_itc_0_clocked_video_vid_f             : out   std_logic;                                        --                                           .vid_f
		vga_alt_vip_itc_0_clocked_video_vid_h             : out   std_logic;                                        --                                           .vid_h
		vga_alt_vip_itc_0_clocked_video_vid_v             : out   std_logic;                                        --                                           .vid_v
		vga_vga_clk_clk                                   : out   std_logic                                         --                                vga_vga_clk.clk
	);
end entity DE1_SoC_QSYS;

architecture rtl of DE1_SoC_QSYS is
	component DE1_SoC_QSYS_audio is
		port (
			clk_clk                      : in  std_logic                     := 'X';             -- clk
			data_divfrec_export          : out std_logic_vector(31 downto 0);                    -- export
			data_fregen_s1_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			data_fregen_s1_write_n       : in  std_logic                     := 'X';             -- write_n
			data_fregen_s1_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			data_fregen_s1_chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_fregen_s1_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			empty_export                 : in  std_logic                     := 'X';             -- export
			empty_s1_address             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			empty_s1_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			fifo_full_export             : in  std_logic                     := 'X';             -- export
			fifo_full_s1_address         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			fifo_full_s1_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			fifo_used_export             : in  std_logic_vector(11 downto 0) := (others => 'X'); -- export
			fifo_used_s1_address         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			fifo_used_s1_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			out_data_audio_export        : out std_logic_vector(31 downto 0);                    -- export
			out_data_audio_s1_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			out_data_audio_s1_write_n    : in  std_logic                     := 'X';             -- write_n
			out_data_audio_s1_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			out_data_audio_s1_chipselect : in  std_logic                     := 'X';             -- chipselect
			out_data_audio_s1_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_pause_export             : out std_logic;                                        -- export
			out_pause_s1_address         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			out_pause_s1_write_n         : in  std_logic                     := 'X';             -- write_n
			out_pause_s1_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			out_pause_s1_chipselect      : in  std_logic                     := 'X';             -- chipselect
			out_pause_s1_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			out_stop_export              : out std_logic;                                        -- export
			out_stop_s1_address          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			out_stop_s1_write_n          : in  std_logic                     := 'X';             -- write_n
			out_stop_s1_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			out_stop_s1_chipselect       : in  std_logic                     := 'X';             -- chipselect
			out_stop_s1_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			reset_reset_n                : in  std_logic                     := 'X';             -- reset_n
			wrclk_export                 : out std_logic;                                        -- export
			wrclk_s1_address             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			wrclk_s1_write_n             : in  std_logic                     := 'X';             -- write_n
			wrclk_s1_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_s1_chipselect          : in  std_logic                     := 'X';             -- chipselect
			wrclk_s1_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			wrreq_export                 : out std_logic;                                        -- export
			wrreq_s1_address             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			wrreq_s1_write_n             : in  std_logic                     := 'X';             -- write_n
			wrreq_s1_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrreq_s1_chipselect          : in  std_logic                     := 'X';             -- chipselect
			wrreq_s1_readdata            : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component DE1_SoC_QSYS_audio;

	component DE1_SoC_QSYS_audio_sel is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component DE1_SoC_QSYS_audio_sel;

	component DE1_SoC_QSYS_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(27 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component DE1_SoC_QSYS_cpu;

	component DE1_SoC_QSYS_dds_increment is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component DE1_SoC_QSYS_dds_increment;

	component DE1_SoC_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_jtag_uart;

	component DE1_SoC_QSYS_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_key;

	component DE1_SoC_QSYS_keyboard_keys is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_keyboard_keys;

	component DE1_SoC_QSYS_lfsr_clk_interrupt_gen is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_lfsr_clk_interrupt_gen;

	component DE1_SoC_QSYS_lfsr_val is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_lfsr_val;

	component DE1_SoC_QSYS_modulation_selector is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component DE1_SoC_QSYS_modulation_selector;

	component DE1_SoC_QSYS_mouse_pos is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_mouse_pos;

	component DE1_SoC_QSYS_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DE1_SoC_QSYS_pll;

	component DE1_SoC_QSYS_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component DE1_SoC_QSYS_sdram;

	component DE1_SoC_QSYS_signal_selector is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component DE1_SoC_QSYS_signal_selector;

	component DE1_SoC_QSYS_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE1_SoC_QSYS_sysid_qsys;

	component DE1_SoC_QSYS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_timer;

	component DE1_SoC_QSYS_vga is
		port (
			alt_vip_itc_0_clocked_video_vid_clk       : in  std_logic                     := 'X';             -- vid_clk
			alt_vip_itc_0_clocked_video_vid_data      : out std_logic_vector(23 downto 0);                    -- vid_data
			alt_vip_itc_0_clocked_video_underflow     : out std_logic;                                        -- underflow
			alt_vip_itc_0_clocked_video_vid_datavalid : out std_logic;                                        -- vid_datavalid
			alt_vip_itc_0_clocked_video_vid_v_sync    : out std_logic;                                        -- vid_v_sync
			alt_vip_itc_0_clocked_video_vid_h_sync    : out std_logic;                                        -- vid_h_sync
			alt_vip_itc_0_clocked_video_vid_f         : out std_logic;                                        -- vid_f
			alt_vip_itc_0_clocked_video_vid_h         : out std_logic;                                        -- vid_h
			alt_vip_itc_0_clocked_video_vid_v         : out std_logic;                                        -- vid_v
			alt_vip_vfr_0_interrupt_sender_irq        : out std_logic;                                        -- irq
			clk_50m_clk                               : in  std_logic                     := 'X';             -- clk
			clk_50m_reset_reset_n                     : in  std_logic                     := 'X';             -- reset_n
			nios_clk_clk                              : in  std_logic                     := 'X';             -- clk
			nios_clk_reset_reset_n                    : in  std_logic                     := 'X';             -- reset_n
			to_nios_2_datamaster_address              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			to_nios_2_datamaster_write                : in  std_logic                     := 'X';             -- write
			to_nios_2_datamaster_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			to_nios_2_datamaster_read                 : in  std_logic                     := 'X';             -- read
			to_nios_2_datamaster_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			to_sdram_address                          : out std_logic_vector(31 downto 0);                    -- address
			to_sdram_burstcount                       : out std_logic_vector(5 downto 0);                     -- burstcount
			to_sdram_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			to_sdram_read                             : out std_logic;                                        -- read
			to_sdram_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			to_sdram_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			vga_clk_clk                               : out std_logic                                         -- clk
		);
	end component DE1_SoC_QSYS_vga;

	component DE1_SoC_QSYS_mm_interconnect_0 is
		port (
			clk_50_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			pll_outclk0_clk                                 : in  std_logic                     := 'X';             -- clk
			pll_outclk2_clk                                 : in  std_logic                     := 'X';             -- clk
			vga_clk_bridge_out_out_clk_1_clk                : in  std_logic                     := 'X';             -- clk
			audio_reset_reset_bridge_in_reset_reset         : in  std_logic                     := 'X';             -- reset
			cpu_reset_n_reset_bridge_in_reset_reset         : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			keyboard_keys_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mouse_pos_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			vga_nios_clk_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                         : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                     : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                            : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                           : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                     : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                  : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest              : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                     : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid            : out std_logic;                                        -- readdatavalid
			vga_to_sdram_address                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vga_to_sdram_waitrequest                        : out std_logic;                                        -- waitrequest
			vga_to_sdram_burstcount                         : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- burstcount
			vga_to_sdram_read                               : in  std_logic                     := 'X';             -- read
			vga_to_sdram_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			vga_to_sdram_readdatavalid                      : out std_logic;                                        -- readdatavalid
			audio_data_fregen_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			audio_data_fregen_s1_write                      : out std_logic;                                        -- write
			audio_data_fregen_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_data_fregen_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			audio_data_fregen_s1_chipselect                 : out std_logic;                                        -- chipselect
			audio_empty_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			audio_empty_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_fifo_full_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			audio_fifo_full_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_fifo_used_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			audio_fifo_used_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_out_data_audio_s1_address                 : out std_logic_vector(1 downto 0);                     -- address
			audio_out_data_audio_s1_write                   : out std_logic;                                        -- write
			audio_out_data_audio_s1_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_out_data_audio_s1_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			audio_out_data_audio_s1_chipselect              : out std_logic;                                        -- chipselect
			audio_out_pause_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			audio_out_pause_s1_write                        : out std_logic;                                        -- write
			audio_out_pause_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_out_pause_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			audio_out_pause_s1_chipselect                   : out std_logic;                                        -- chipselect
			audio_out_stop_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			audio_out_stop_s1_write                         : out std_logic;                                        -- write
			audio_out_stop_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_out_stop_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			audio_out_stop_s1_chipselect                    : out std_logic;                                        -- chipselect
			audio_wrclk_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			audio_wrclk_s1_write                            : out std_logic;                                        -- write
			audio_wrclk_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_wrclk_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			audio_wrclk_s1_chipselect                       : out std_logic;                                        -- chipselect
			audio_wrreq_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			audio_wrreq_s1_write                            : out std_logic;                                        -- write
			audio_wrreq_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_wrreq_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			audio_wrreq_s1_chipselect                       : out std_logic;                                        -- chipselect
			audio_sel_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			audio_sel_s1_write                              : out std_logic;                                        -- write
			audio_sel_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_sel_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			audio_sel_s1_chipselect                         : out std_logic;                                        -- chipselect
			cpu_jtag_debug_module_address                   : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write                     : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                      : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess               : out std_logic;                                        -- debugaccess
			dds_increment_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			dds_increment_s1_write                          : out std_logic;                                        -- write
			dds_increment_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dds_increment_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			dds_increment_s1_chipselect                     : out std_logic;                                        -- chipselect
			div_freq_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			div_freq_s1_write                               : out std_logic;                                        -- write
			div_freq_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			div_freq_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			div_freq_s1_chipselect                          : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write               : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			key_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                    : out std_logic;                                        -- write
			key_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                               : out std_logic;                                        -- chipselect
			keyboard_keys_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			keyboard_keys_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lfsr_clk_interrupt_gen_s1_address               : out std_logic_vector(1 downto 0);                     -- address
			lfsr_clk_interrupt_gen_s1_write                 : out std_logic;                                        -- write
			lfsr_clk_interrupt_gen_s1_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lfsr_clk_interrupt_gen_s1_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			lfsr_clk_interrupt_gen_s1_chipselect            : out std_logic;                                        -- chipselect
			lfsr_val_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			lfsr_val_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			modulation_selector_s1_address                  : out std_logic_vector(1 downto 0);                     -- address
			modulation_selector_s1_write                    : out std_logic;                                        -- write
			modulation_selector_s1_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			modulation_selector_s1_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			modulation_selector_s1_chipselect               : out std_logic;                                        -- chipselect
			mouse_pos_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			mouse_pos_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_address                                : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                  : out std_logic;                                        -- write
			sdram_s1_read                                   : out std_logic;                                        -- read
			sdram_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                             : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                             : out std_logic;                                        -- chipselect
			signal_selector_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			signal_selector_s1_write                        : out std_logic;                                        -- write
			signal_selector_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			signal_selector_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			signal_selector_s1_chipselect                   : out std_logic;                                        -- chipselect
			sysid_qsys_control_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                                : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                  : out std_logic;                                        -- write
			timer_s1_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                             : out std_logic;                                        -- chipselect
			vga_to_nios_2_datamaster_address                : out std_logic_vector(4 downto 0);                     -- address
			vga_to_nios_2_datamaster_write                  : out std_logic;                                        -- write
			vga_to_nios_2_datamaster_read                   : out std_logic;                                        -- read
			vga_to_nios_2_datamaster_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vga_to_nios_2_datamaster_writedata              : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component DE1_SoC_QSYS_mm_interconnect_0;

	component DE1_SoC_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE1_SoC_QSYS_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component de1_soc_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de1_soc_qsys_rst_controller;

	component de1_soc_qsys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de1_soc_qsys_rst_controller_002;

	signal pll_outclk0_clk                                               : std_logic;                     -- pll:outclk_0 -> [audio:clk_clk, irq_synchronizer:receiver_clk, mm_interconnect_0:pll_outclk0_clk, rst_controller:clk, sdram:clk, vga:nios_clk_clk]
	signal pll_outclk2_clk                                               : std_logic;                     -- pll:outclk_2 -> [clk_25_out_clk, keyboard_keys:clk, mm_interconnect_0:pll_outclk2_clk, rst_controller_003:clk]
	signal vga_vga_clk_clk_internal                                      : std_logic;                     -- vga:vga_clk_clk -> [vga_vga_clk_clk, mm_interconnect_0:vga_clk_bridge_out_out_clk_1_clk, mouse_pos:clk, rst_controller_004:clk]
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal vga_to_sdram_readdata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_to_sdram_readdata -> vga:to_sdram_readdata
	signal vga_to_sdram_waitrequest                                      : std_logic;                     -- mm_interconnect_0:vga_to_sdram_waitrequest -> vga:to_sdram_waitrequest
	signal vga_to_sdram_address                                          : std_logic_vector(31 downto 0); -- vga:to_sdram_address -> mm_interconnect_0:vga_to_sdram_address
	signal vga_to_sdram_read                                             : std_logic;                     -- vga:to_sdram_read -> mm_interconnect_0:vga_to_sdram_read
	signal vga_to_sdram_readdatavalid                                    : std_logic;                     -- mm_interconnect_0:vga_to_sdram_readdatavalid -> vga:to_sdram_readdatavalid
	signal vga_to_sdram_burstcount                                       : std_logic_vector(5 downto 0);  -- vga:to_sdram_burstcount -> mm_interconnect_0:vga_to_sdram_burstcount
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_audio_data_fregen_s1_chipselect             : std_logic;                     -- mm_interconnect_0:audio_data_fregen_s1_chipselect -> audio:data_fregen_s1_chipselect
	signal mm_interconnect_0_audio_data_fregen_s1_readdata               : std_logic_vector(31 downto 0); -- audio:data_fregen_s1_readdata -> mm_interconnect_0:audio_data_fregen_s1_readdata
	signal mm_interconnect_0_audio_data_fregen_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_data_fregen_s1_address -> audio:data_fregen_s1_address
	signal mm_interconnect_0_audio_data_fregen_s1_write                  : std_logic;                     -- mm_interconnect_0:audio_data_fregen_s1_write -> mm_interconnect_0_audio_data_fregen_s1_write:in
	signal mm_interconnect_0_audio_data_fregen_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_data_fregen_s1_writedata -> audio:data_fregen_s1_writedata
	signal mm_interconnect_0_audio_empty_s1_readdata                     : std_logic_vector(31 downto 0); -- audio:empty_s1_readdata -> mm_interconnect_0:audio_empty_s1_readdata
	signal mm_interconnect_0_audio_empty_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_empty_s1_address -> audio:empty_s1_address
	signal mm_interconnect_0_audio_fifo_full_s1_readdata                 : std_logic_vector(31 downto 0); -- audio:fifo_full_s1_readdata -> mm_interconnect_0:audio_fifo_full_s1_readdata
	signal mm_interconnect_0_audio_fifo_full_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_fifo_full_s1_address -> audio:fifo_full_s1_address
	signal mm_interconnect_0_audio_fifo_used_s1_readdata                 : std_logic_vector(31 downto 0); -- audio:fifo_used_s1_readdata -> mm_interconnect_0:audio_fifo_used_s1_readdata
	signal mm_interconnect_0_audio_fifo_used_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_fifo_used_s1_address -> audio:fifo_used_s1_address
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata              : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest           : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess           : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_read                  : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_0_cpu_jtag_debug_module_write                 : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_0_audio_out_data_audio_s1_chipselect          : std_logic;                     -- mm_interconnect_0:audio_out_data_audio_s1_chipselect -> audio:out_data_audio_s1_chipselect
	signal mm_interconnect_0_audio_out_data_audio_s1_readdata            : std_logic_vector(31 downto 0); -- audio:out_data_audio_s1_readdata -> mm_interconnect_0:audio_out_data_audio_s1_readdata
	signal mm_interconnect_0_audio_out_data_audio_s1_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_out_data_audio_s1_address -> audio:out_data_audio_s1_address
	signal mm_interconnect_0_audio_out_data_audio_s1_write               : std_logic;                     -- mm_interconnect_0:audio_out_data_audio_s1_write -> mm_interconnect_0_audio_out_data_audio_s1_write:in
	signal mm_interconnect_0_audio_out_data_audio_s1_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_out_data_audio_s1_writedata -> audio:out_data_audio_s1_writedata
	signal mm_interconnect_0_audio_out_pause_s1_chipselect               : std_logic;                     -- mm_interconnect_0:audio_out_pause_s1_chipselect -> audio:out_pause_s1_chipselect
	signal mm_interconnect_0_audio_out_pause_s1_readdata                 : std_logic_vector(31 downto 0); -- audio:out_pause_s1_readdata -> mm_interconnect_0:audio_out_pause_s1_readdata
	signal mm_interconnect_0_audio_out_pause_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_out_pause_s1_address -> audio:out_pause_s1_address
	signal mm_interconnect_0_audio_out_pause_s1_write                    : std_logic;                     -- mm_interconnect_0:audio_out_pause_s1_write -> mm_interconnect_0_audio_out_pause_s1_write:in
	signal mm_interconnect_0_audio_out_pause_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_out_pause_s1_writedata -> audio:out_pause_s1_writedata
	signal mm_interconnect_0_audio_out_stop_s1_chipselect                : std_logic;                     -- mm_interconnect_0:audio_out_stop_s1_chipselect -> audio:out_stop_s1_chipselect
	signal mm_interconnect_0_audio_out_stop_s1_readdata                  : std_logic_vector(31 downto 0); -- audio:out_stop_s1_readdata -> mm_interconnect_0:audio_out_stop_s1_readdata
	signal mm_interconnect_0_audio_out_stop_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_out_stop_s1_address -> audio:out_stop_s1_address
	signal mm_interconnect_0_audio_out_stop_s1_write                     : std_logic;                     -- mm_interconnect_0:audio_out_stop_s1_write -> mm_interconnect_0_audio_out_stop_s1_write:in
	signal mm_interconnect_0_audio_out_stop_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_out_stop_s1_writedata -> audio:out_stop_s1_writedata
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_0_key_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                             : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_signal_selector_s1_chipselect               : std_logic;                     -- mm_interconnect_0:signal_selector_s1_chipselect -> signal_selector:chipselect
	signal mm_interconnect_0_signal_selector_s1_readdata                 : std_logic_vector(31 downto 0); -- signal_selector:readdata -> mm_interconnect_0:signal_selector_s1_readdata
	signal mm_interconnect_0_signal_selector_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:signal_selector_s1_address -> signal_selector:address
	signal mm_interconnect_0_signal_selector_s1_write                    : std_logic;                     -- mm_interconnect_0:signal_selector_s1_write -> mm_interconnect_0_signal_selector_s1_write:in
	signal mm_interconnect_0_signal_selector_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:signal_selector_s1_writedata -> signal_selector:writedata
	signal mm_interconnect_0_modulation_selector_s1_chipselect           : std_logic;                     -- mm_interconnect_0:modulation_selector_s1_chipselect -> modulation_selector:chipselect
	signal mm_interconnect_0_modulation_selector_s1_readdata             : std_logic_vector(31 downto 0); -- modulation_selector:readdata -> mm_interconnect_0:modulation_selector_s1_readdata
	signal mm_interconnect_0_modulation_selector_s1_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:modulation_selector_s1_address -> modulation_selector:address
	signal mm_interconnect_0_modulation_selector_s1_write                : std_logic;                     -- mm_interconnect_0:modulation_selector_s1_write -> mm_interconnect_0_modulation_selector_s1_write:in
	signal mm_interconnect_0_modulation_selector_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:modulation_selector_s1_writedata -> modulation_selector:writedata
	signal mm_interconnect_0_keyboard_keys_s1_readdata                   : std_logic_vector(31 downto 0); -- keyboard_keys:readdata -> mm_interconnect_0:keyboard_keys_s1_readdata
	signal mm_interconnect_0_keyboard_keys_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:keyboard_keys_s1_address -> keyboard_keys:address
	signal mm_interconnect_0_mouse_pos_s1_readdata                       : std_logic_vector(31 downto 0); -- mouse_pos:readdata -> mm_interconnect_0:mouse_pos_s1_readdata
	signal mm_interconnect_0_mouse_pos_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:mouse_pos_s1_address -> mouse_pos:address
	signal mm_interconnect_0_div_freq_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:div_freq_s1_chipselect -> div_freq:chipselect
	signal mm_interconnect_0_div_freq_s1_readdata                        : std_logic_vector(31 downto 0); -- div_freq:readdata -> mm_interconnect_0:div_freq_s1_readdata
	signal mm_interconnect_0_div_freq_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:div_freq_s1_address -> div_freq:address
	signal mm_interconnect_0_div_freq_s1_write                           : std_logic;                     -- mm_interconnect_0:div_freq_s1_write -> mm_interconnect_0_div_freq_s1_write:in
	signal mm_interconnect_0_div_freq_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:div_freq_s1_writedata -> div_freq:writedata
	signal mm_interconnect_0_audio_sel_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:audio_sel_s1_chipselect -> audio_sel:chipselect
	signal mm_interconnect_0_audio_sel_s1_readdata                       : std_logic_vector(31 downto 0); -- audio_sel:readdata -> mm_interconnect_0:audio_sel_s1_readdata
	signal mm_interconnect_0_audio_sel_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_sel_s1_address -> audio_sel:address
	signal mm_interconnect_0_audio_sel_s1_write                          : std_logic;                     -- mm_interconnect_0:audio_sel_s1_write -> mm_interconnect_0_audio_sel_s1_write:in
	signal mm_interconnect_0_audio_sel_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_sel_s1_writedata -> audio_sel:writedata
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect        : std_logic;                     -- mm_interconnect_0:lfsr_clk_interrupt_gen_s1_chipselect -> lfsr_clk_interrupt_gen:chipselect
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata          : std_logic_vector(31 downto 0); -- lfsr_clk_interrupt_gen:readdata -> mm_interconnect_0:lfsr_clk_interrupt_gen_s1_readdata
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:lfsr_clk_interrupt_gen_s1_address -> lfsr_clk_interrupt_gen:address
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write             : std_logic;                     -- mm_interconnect_0:lfsr_clk_interrupt_gen_s1_write -> mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write:in
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:lfsr_clk_interrupt_gen_s1_writedata -> lfsr_clk_interrupt_gen:writedata
	signal mm_interconnect_0_lfsr_val_s1_readdata                        : std_logic_vector(31 downto 0); -- lfsr_val:readdata -> mm_interconnect_0:lfsr_val_s1_readdata
	signal mm_interconnect_0_lfsr_val_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:lfsr_val_s1_address -> lfsr_val:address
	signal mm_interconnect_0_dds_increment_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:dds_increment_s1_chipselect -> dds_increment:chipselect
	signal mm_interconnect_0_dds_increment_s1_readdata                   : std_logic_vector(31 downto 0); -- dds_increment:readdata -> mm_interconnect_0:dds_increment_s1_readdata
	signal mm_interconnect_0_dds_increment_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:dds_increment_s1_address -> dds_increment:address
	signal mm_interconnect_0_dds_increment_s1_write                      : std_logic;                     -- mm_interconnect_0:dds_increment_s1_write -> mm_interconnect_0_dds_increment_s1_write:in
	signal mm_interconnect_0_dds_increment_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:dds_increment_s1_writedata -> dds_increment:writedata
	signal mm_interconnect_0_vga_to_nios_2_datamaster_readdata           : std_logic_vector(31 downto 0); -- vga:to_nios_2_datamaster_readdata -> mm_interconnect_0:vga_to_nios_2_datamaster_readdata
	signal mm_interconnect_0_vga_to_nios_2_datamaster_address            : std_logic_vector(4 downto 0);  -- mm_interconnect_0:vga_to_nios_2_datamaster_address -> vga:to_nios_2_datamaster_address
	signal mm_interconnect_0_vga_to_nios_2_datamaster_read               : std_logic;                     -- mm_interconnect_0:vga_to_nios_2_datamaster_read -> vga:to_nios_2_datamaster_read
	signal mm_interconnect_0_vga_to_nios_2_datamaster_write              : std_logic;                     -- mm_interconnect_0:vga_to_nios_2_datamaster_write -> vga:to_nios_2_datamaster_write
	signal mm_interconnect_0_vga_to_nios_2_datamaster_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:vga_to_nios_2_datamaster_writedata -> vga:to_nios_2_datamaster_writedata
	signal mm_interconnect_0_audio_wrclk_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:audio_wrclk_s1_chipselect -> audio:wrclk_s1_chipselect
	signal mm_interconnect_0_audio_wrclk_s1_readdata                     : std_logic_vector(31 downto 0); -- audio:wrclk_s1_readdata -> mm_interconnect_0:audio_wrclk_s1_readdata
	signal mm_interconnect_0_audio_wrclk_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_wrclk_s1_address -> audio:wrclk_s1_address
	signal mm_interconnect_0_audio_wrclk_s1_write                        : std_logic;                     -- mm_interconnect_0:audio_wrclk_s1_write -> mm_interconnect_0_audio_wrclk_s1_write:in
	signal mm_interconnect_0_audio_wrclk_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_wrclk_s1_writedata -> audio:wrclk_s1_writedata
	signal mm_interconnect_0_audio_wrreq_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:audio_wrreq_s1_chipselect -> audio:wrreq_s1_chipselect
	signal mm_interconnect_0_audio_wrreq_s1_readdata                     : std_logic_vector(31 downto 0); -- audio:wrreq_s1_readdata -> mm_interconnect_0:audio_wrreq_s1_readdata
	signal mm_interconnect_0_audio_wrreq_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_wrreq_s1_address -> audio:wrreq_s1_address
	signal mm_interconnect_0_audio_wrreq_s1_write                        : std_logic;                     -- mm_interconnect_0:audio_wrreq_s1_write -> mm_interconnect_0_audio_wrreq_s1_write:in
	signal mm_interconnect_0_audio_wrreq_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_wrreq_s1_writedata -> audio:wrreq_s1_writedata
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- key:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                      : std_logic;                     -- lfsr_clk_interrupt_gen:irq -> irq_mapper:receiver4_irq
	signal cpu_d_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                 : std_logic_vector(0 downto 0);  -- vga:alt_vip_vfr_0_interrupt_sender_irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:audio_reset_reset_bridge_in_reset_reset, mm_interconnect_0:vga_nios_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                            : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_002_reset_out_reset_req                        : std_logic;                     -- rst_controller_002:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal cpu_jtag_debug_module_reset_reset                             : std_logic;                     -- cpu:jtag_debug_module_resetrequest -> rst_controller_002:reset_in1
	signal rst_controller_003_reset_out_reset                            : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:keyboard_keys_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal rst_controller_004_reset_out_reset                            : std_logic;                     -- rst_controller_004:reset_out -> [mm_interconnect_0:mouse_pos_reset_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_audio_data_fregen_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_audio_data_fregen_s1_write:inv -> audio:data_fregen_s1_write_n
	signal mm_interconnect_0_audio_out_data_audio_s1_write_ports_inv     : std_logic;                     -- mm_interconnect_0_audio_out_data_audio_s1_write:inv -> audio:out_data_audio_s1_write_n
	signal mm_interconnect_0_audio_out_pause_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_audio_out_pause_s1_write:inv -> audio:out_pause_s1_write_n
	signal mm_interconnect_0_audio_out_stop_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_audio_out_stop_s1_write:inv -> audio:out_stop_s1_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_signal_selector_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_signal_selector_s1_write:inv -> signal_selector:write_n
	signal mm_interconnect_0_modulation_selector_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_modulation_selector_s1_write:inv -> modulation_selector:write_n
	signal mm_interconnect_0_div_freq_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_div_freq_s1_write:inv -> div_freq:write_n
	signal mm_interconnect_0_audio_sel_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_audio_sel_s1_write:inv -> audio_sel:write_n
	signal mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write:inv -> lfsr_clk_interrupt_gen:write_n
	signal mm_interconnect_0_dds_increment_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_dds_increment_s1_write:inv -> dds_increment:write_n
	signal mm_interconnect_0_audio_wrclk_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_audio_wrclk_s1_write:inv -> audio:wrclk_s1_write_n
	signal mm_interconnect_0_audio_wrreq_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_audio_wrreq_s1_write:inv -> audio:wrreq_s1_write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [audio:reset_reset_n, sdram:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [audio_sel:reset_n, dds_increment:reset_n, div_freq:reset_n, jtag_uart:rst_n, key:reset_n, lfsr_clk_interrupt_gen:reset_n, lfsr_val:reset_n, modulation_selector:reset_n, signal_selector:reset_n, sysid_qsys:reset_n, timer:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> cpu:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> keyboard_keys:reset_n
	signal rst_controller_004_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> mouse_pos:reset_n

begin

	audio : component DE1_SoC_QSYS_audio
		port map (
			clk_clk                      => pll_outclk0_clk,                                           --               clk.clk
			data_divfrec_export          => audio2fifo_0_data_divfrec_export,                          --      data_divfrec.export
			data_fregen_s1_address       => mm_interconnect_0_audio_data_fregen_s1_address,            --    data_fregen_s1.address
			data_fregen_s1_write_n       => mm_interconnect_0_audio_data_fregen_s1_write_ports_inv,    --                  .write_n
			data_fregen_s1_writedata     => mm_interconnect_0_audio_data_fregen_s1_writedata,          --                  .writedata
			data_fregen_s1_chipselect    => mm_interconnect_0_audio_data_fregen_s1_chipselect,         --                  .chipselect
			data_fregen_s1_readdata      => mm_interconnect_0_audio_data_fregen_s1_readdata,           --                  .readdata
			empty_export                 => audio2fifo_0_empty_export,                                 --             empty.export
			empty_s1_address             => mm_interconnect_0_audio_empty_s1_address,                  --          empty_s1.address
			empty_s1_readdata            => mm_interconnect_0_audio_empty_s1_readdata,                 --                  .readdata
			fifo_full_export             => audio2fifo_0_fifo_full_export,                             --         fifo_full.export
			fifo_full_s1_address         => mm_interconnect_0_audio_fifo_full_s1_address,              --      fifo_full_s1.address
			fifo_full_s1_readdata        => mm_interconnect_0_audio_fifo_full_s1_readdata,             --                  .readdata
			fifo_used_export             => audio2fifo_0_fifo_used_export,                             --         fifo_used.export
			fifo_used_s1_address         => mm_interconnect_0_audio_fifo_used_s1_address,              --      fifo_used_s1.address
			fifo_used_s1_readdata        => mm_interconnect_0_audio_fifo_used_s1_readdata,             --                  .readdata
			out_data_audio_export        => audio2fifo_0_out_data_audio_export,                        --    out_data_audio.export
			out_data_audio_s1_address    => mm_interconnect_0_audio_out_data_audio_s1_address,         -- out_data_audio_s1.address
			out_data_audio_s1_write_n    => mm_interconnect_0_audio_out_data_audio_s1_write_ports_inv, --                  .write_n
			out_data_audio_s1_writedata  => mm_interconnect_0_audio_out_data_audio_s1_writedata,       --                  .writedata
			out_data_audio_s1_chipselect => mm_interconnect_0_audio_out_data_audio_s1_chipselect,      --                  .chipselect
			out_data_audio_s1_readdata   => mm_interconnect_0_audio_out_data_audio_s1_readdata,        --                  .readdata
			out_pause_export             => audio2fifo_0_out_pause_export,                             --         out_pause.export
			out_pause_s1_address         => mm_interconnect_0_audio_out_pause_s1_address,              --      out_pause_s1.address
			out_pause_s1_write_n         => mm_interconnect_0_audio_out_pause_s1_write_ports_inv,      --                  .write_n
			out_pause_s1_writedata       => mm_interconnect_0_audio_out_pause_s1_writedata,            --                  .writedata
			out_pause_s1_chipselect      => mm_interconnect_0_audio_out_pause_s1_chipselect,           --                  .chipselect
			out_pause_s1_readdata        => mm_interconnect_0_audio_out_pause_s1_readdata,             --                  .readdata
			out_stop_export              => audio2fifo_0_out_stop_export,                              --          out_stop.export
			out_stop_s1_address          => mm_interconnect_0_audio_out_stop_s1_address,               --       out_stop_s1.address
			out_stop_s1_write_n          => mm_interconnect_0_audio_out_stop_s1_write_ports_inv,       --                  .write_n
			out_stop_s1_writedata        => mm_interconnect_0_audio_out_stop_s1_writedata,             --                  .writedata
			out_stop_s1_chipselect       => mm_interconnect_0_audio_out_stop_s1_chipselect,            --                  .chipselect
			out_stop_s1_readdata         => mm_interconnect_0_audio_out_stop_s1_readdata,              --                  .readdata
			reset_reset_n                => rst_controller_reset_out_reset_ports_inv,                  --             reset.reset_n
			wrclk_export                 => audio2fifo_0_wrclk_export,                                 --             wrclk.export
			wrclk_s1_address             => mm_interconnect_0_audio_wrclk_s1_address,                  --          wrclk_s1.address
			wrclk_s1_write_n             => mm_interconnect_0_audio_wrclk_s1_write_ports_inv,          --                  .write_n
			wrclk_s1_writedata           => mm_interconnect_0_audio_wrclk_s1_writedata,                --                  .writedata
			wrclk_s1_chipselect          => mm_interconnect_0_audio_wrclk_s1_chipselect,               --                  .chipselect
			wrclk_s1_readdata            => mm_interconnect_0_audio_wrclk_s1_readdata,                 --                  .readdata
			wrreq_export                 => audio2fifo_0_wrreq_export,                                 --             wrreq.export
			wrreq_s1_address             => mm_interconnect_0_audio_wrreq_s1_address,                  --          wrreq_s1.address
			wrreq_s1_write_n             => mm_interconnect_0_audio_wrreq_s1_write_ports_inv,          --                  .write_n
			wrreq_s1_writedata           => mm_interconnect_0_audio_wrreq_s1_writedata,                --                  .writedata
			wrreq_s1_chipselect          => mm_interconnect_0_audio_wrreq_s1_chipselect,               --                  .chipselect
			wrreq_s1_readdata            => mm_interconnect_0_audio_wrreq_s1_readdata                  --                  .readdata
		);

	audio_sel : component DE1_SoC_QSYS_audio_sel
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_audio_sel_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_audio_sel_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_audio_sel_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_audio_sel_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_audio_sel_s1_readdata,        --                    .readdata
			out_port   => audio_sel_export                                -- external_connection.export
		);

	cpu : component DE1_SoC_QSYS_cpu
		port map (
			clk                                   => clk_clk,                                             --                       clk.clk
			reset_n                               => rst_controller_002_reset_out_reset_ports_inv,        --                   reset_n.reset_n
			reset_req                             => rst_controller_002_reset_out_reset_req,              --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			d_readdatavalid                       => cpu_data_master_readdatavalid,                       --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	dds_increment : component DE1_SoC_QSYS_dds_increment
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_dds_increment_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_dds_increment_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_dds_increment_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_dds_increment_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_dds_increment_s1_readdata,        --                    .readdata
			out_port   => dds_increment_external_connection_export            -- external_connection.export
		);

	div_freq : component DE1_SoC_QSYS_dds_increment
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_div_freq_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_div_freq_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_div_freq_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_div_freq_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_div_freq_s1_readdata,        --                    .readdata
			out_port   => div_freq_export                                -- external_connection.export
		);

	jtag_uart : component DE1_SoC_QSYS_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	key : component DE1_SoC_QSYS_key
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,             --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,            --                    .readdata
			in_port    => key_external_connection_export,               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	keyboard_keys : component DE1_SoC_QSYS_keyboard_keys
		port map (
			clk      => pll_outclk2_clk,                              --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_keyboard_keys_s1_address,   --                  s1.address
			readdata => mm_interconnect_0_keyboard_keys_s1_readdata,  --                    .readdata
			in_port  => keyboard_keys_export                          -- external_connection.export
		);

	lfsr_clk_interrupt_gen : component DE1_SoC_QSYS_lfsr_clk_interrupt_gen
		port map (
			clk        => clk_clk,                                                     --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata,        --                    .readdata
			in_port    => lfsr_clk_interrupt_gen_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver4_irq                                     --                 irq.irq
		);

	lfsr_val : component DE1_SoC_QSYS_lfsr_val
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_lfsr_val_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_lfsr_val_s1_readdata,       --                    .readdata
			in_port  => lfsr_val_external_connection_export           -- external_connection.export
		);

	modulation_selector : component DE1_SoC_QSYS_modulation_selector
		port map (
			clk        => clk_clk,                                                  --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_modulation_selector_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_modulation_selector_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_modulation_selector_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_modulation_selector_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_modulation_selector_s1_readdata,        --                    .readdata
			out_port   => modulation_selector_export                                -- external_connection.export
		);

	mouse_pos : component DE1_SoC_QSYS_mouse_pos
		port map (
			clk      => vga_vga_clk_clk_internal,                     --                 clk.clk
			reset_n  => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_mouse_pos_s1_address,       --                  s1.address
			readdata => mm_interconnect_0_mouse_pos_s1_readdata,      --                    .readdata
			in_port  => mouse_pos_export                              -- external_connection.export
		);

	pll : component DE1_SoC_QSYS_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => clk_sdram_clk,           -- outclk1.clk
			outclk_2 => pll_outclk2_clk,         -- outclk2.clk
			locked   => pll_locked_export        --  locked.export
		);

	sdram : component DE1_SoC_QSYS_sdram
		port map (
			clk            => pll_outclk0_clk,                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	signal_selector : component DE1_SoC_QSYS_signal_selector
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_signal_selector_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_signal_selector_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_signal_selector_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_signal_selector_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_signal_selector_s1_readdata,        --                    .readdata
			out_port   => signal_selector_export                                -- external_connection.export
		);

	sysid_qsys : component DE1_SoC_QSYS_sysid_qsys
		port map (
			clock    => clk_clk,                                               --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer : component DE1_SoC_QSYS_timer
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,           --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,         --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,          --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,        --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv,   --      .write_n
			irq        => irq_mapper_receiver2_irq                      --   irq.irq
		);

	vga : component DE1_SoC_QSYS_vga
		port map (
			alt_vip_itc_0_clocked_video_vid_clk       => vga_alt_vip_itc_0_clocked_video_vid_clk,              --    alt_vip_itc_0_clocked_video.vid_clk
			alt_vip_itc_0_clocked_video_vid_data      => vga_alt_vip_itc_0_clocked_video_vid_data,             --                               .vid_data
			alt_vip_itc_0_clocked_video_underflow     => vga_alt_vip_itc_0_clocked_video_underflow,            --                               .underflow
			alt_vip_itc_0_clocked_video_vid_datavalid => vga_alt_vip_itc_0_clocked_video_vid_datavalid,        --                               .vid_datavalid
			alt_vip_itc_0_clocked_video_vid_v_sync    => vga_alt_vip_itc_0_clocked_video_vid_v_sync,           --                               .vid_v_sync
			alt_vip_itc_0_clocked_video_vid_h_sync    => vga_alt_vip_itc_0_clocked_video_vid_h_sync,           --                               .vid_h_sync
			alt_vip_itc_0_clocked_video_vid_f         => vga_alt_vip_itc_0_clocked_video_vid_f,                --                               .vid_f
			alt_vip_itc_0_clocked_video_vid_h         => vga_alt_vip_itc_0_clocked_video_vid_h,                --                               .vid_h
			alt_vip_itc_0_clocked_video_vid_v         => vga_alt_vip_itc_0_clocked_video_vid_v,                --                               .vid_v
			alt_vip_vfr_0_interrupt_sender_irq        => irq_synchronizer_receiver_irq(0),                     -- alt_vip_vfr_0_interrupt_sender.irq
			clk_50m_clk                               => clk_clk,                                              --                        clk_50m.clk
			clk_50m_reset_reset_n                     => reset_reset_n,                                        --                  clk_50m_reset.reset_n
			nios_clk_clk                              => pll_outclk0_clk,                                      --                       nios_clk.clk
			nios_clk_reset_reset_n                    => reset_reset_n,                                        --                 nios_clk_reset.reset_n
			to_nios_2_datamaster_address              => mm_interconnect_0_vga_to_nios_2_datamaster_address,   --           to_nios_2_datamaster.address
			to_nios_2_datamaster_write                => mm_interconnect_0_vga_to_nios_2_datamaster_write,     --                               .write
			to_nios_2_datamaster_writedata            => mm_interconnect_0_vga_to_nios_2_datamaster_writedata, --                               .writedata
			to_nios_2_datamaster_read                 => mm_interconnect_0_vga_to_nios_2_datamaster_read,      --                               .read
			to_nios_2_datamaster_readdata             => mm_interconnect_0_vga_to_nios_2_datamaster_readdata,  --                               .readdata
			to_sdram_address                          => vga_to_sdram_address,                                 --                       to_sdram.address
			to_sdram_burstcount                       => vga_to_sdram_burstcount,                              --                               .burstcount
			to_sdram_readdata                         => vga_to_sdram_readdata,                                --                               .readdata
			to_sdram_read                             => vga_to_sdram_read,                                    --                               .read
			to_sdram_readdatavalid                    => vga_to_sdram_readdatavalid,                           --                               .readdatavalid
			to_sdram_waitrequest                      => vga_to_sdram_waitrequest,                             --                               .waitrequest
			vga_clk_clk                               => vga_vga_clk_clk_internal                              --                        vga_clk.clk
		);

	mm_interconnect_0 : component DE1_SoC_QSYS_mm_interconnect_0
		port map (
			clk_50_clk_clk                                  => clk_clk,                                                   --                                clk_50_clk.clk
			pll_outclk0_clk                                 => pll_outclk0_clk,                                           --                               pll_outclk0.clk
			pll_outclk2_clk                                 => pll_outclk2_clk,                                           --                               pll_outclk2.clk
			vga_clk_bridge_out_out_clk_1_clk                => vga_vga_clk_clk_internal,                                  --              vga_clk_bridge_out_out_clk_1.clk
			audio_reset_reset_bridge_in_reset_reset         => rst_controller_reset_out_reset,                            --         audio_reset_reset_bridge_in_reset.reset
			cpu_reset_n_reset_bridge_in_reset_reset         => rst_controller_002_reset_out_reset,                        --         cpu_reset_n_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset     => rst_controller_001_reset_out_reset,                        --     jtag_uart_reset_reset_bridge_in_reset.reset
			keyboard_keys_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                        -- keyboard_keys_reset_reset_bridge_in_reset.reset
			mouse_pos_reset_reset_bridge_in_reset_reset     => rst_controller_004_reset_out_reset,                        --     mouse_pos_reset_reset_bridge_in_reset.reset
			vga_nios_clk_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                            --  vga_nios_clk_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                         => cpu_data_master_address,                                   --                           cpu_data_master.address
			cpu_data_master_waitrequest                     => cpu_data_master_waitrequest,                               --                                          .waitrequest
			cpu_data_master_byteenable                      => cpu_data_master_byteenable,                                --                                          .byteenable
			cpu_data_master_read                            => cpu_data_master_read,                                      --                                          .read
			cpu_data_master_readdata                        => cpu_data_master_readdata,                                  --                                          .readdata
			cpu_data_master_readdatavalid                   => cpu_data_master_readdatavalid,                             --                                          .readdatavalid
			cpu_data_master_write                           => cpu_data_master_write,                                     --                                          .write
			cpu_data_master_writedata                       => cpu_data_master_writedata,                                 --                                          .writedata
			cpu_data_master_debugaccess                     => cpu_data_master_debugaccess,                               --                                          .debugaccess
			cpu_instruction_master_address                  => cpu_instruction_master_address,                            --                    cpu_instruction_master.address
			cpu_instruction_master_waitrequest              => cpu_instruction_master_waitrequest,                        --                                          .waitrequest
			cpu_instruction_master_read                     => cpu_instruction_master_read,                               --                                          .read
			cpu_instruction_master_readdata                 => cpu_instruction_master_readdata,                           --                                          .readdata
			cpu_instruction_master_readdatavalid            => cpu_instruction_master_readdatavalid,                      --                                          .readdatavalid
			vga_to_sdram_address                            => vga_to_sdram_address,                                      --                              vga_to_sdram.address
			vga_to_sdram_waitrequest                        => vga_to_sdram_waitrequest,                                  --                                          .waitrequest
			vga_to_sdram_burstcount                         => vga_to_sdram_burstcount,                                   --                                          .burstcount
			vga_to_sdram_read                               => vga_to_sdram_read,                                         --                                          .read
			vga_to_sdram_readdata                           => vga_to_sdram_readdata,                                     --                                          .readdata
			vga_to_sdram_readdatavalid                      => vga_to_sdram_readdatavalid,                                --                                          .readdatavalid
			audio_data_fregen_s1_address                    => mm_interconnect_0_audio_data_fregen_s1_address,            --                      audio_data_fregen_s1.address
			audio_data_fregen_s1_write                      => mm_interconnect_0_audio_data_fregen_s1_write,              --                                          .write
			audio_data_fregen_s1_readdata                   => mm_interconnect_0_audio_data_fregen_s1_readdata,           --                                          .readdata
			audio_data_fregen_s1_writedata                  => mm_interconnect_0_audio_data_fregen_s1_writedata,          --                                          .writedata
			audio_data_fregen_s1_chipselect                 => mm_interconnect_0_audio_data_fregen_s1_chipselect,         --                                          .chipselect
			audio_empty_s1_address                          => mm_interconnect_0_audio_empty_s1_address,                  --                            audio_empty_s1.address
			audio_empty_s1_readdata                         => mm_interconnect_0_audio_empty_s1_readdata,                 --                                          .readdata
			audio_fifo_full_s1_address                      => mm_interconnect_0_audio_fifo_full_s1_address,              --                        audio_fifo_full_s1.address
			audio_fifo_full_s1_readdata                     => mm_interconnect_0_audio_fifo_full_s1_readdata,             --                                          .readdata
			audio_fifo_used_s1_address                      => mm_interconnect_0_audio_fifo_used_s1_address,              --                        audio_fifo_used_s1.address
			audio_fifo_used_s1_readdata                     => mm_interconnect_0_audio_fifo_used_s1_readdata,             --                                          .readdata
			audio_out_data_audio_s1_address                 => mm_interconnect_0_audio_out_data_audio_s1_address,         --                   audio_out_data_audio_s1.address
			audio_out_data_audio_s1_write                   => mm_interconnect_0_audio_out_data_audio_s1_write,           --                                          .write
			audio_out_data_audio_s1_readdata                => mm_interconnect_0_audio_out_data_audio_s1_readdata,        --                                          .readdata
			audio_out_data_audio_s1_writedata               => mm_interconnect_0_audio_out_data_audio_s1_writedata,       --                                          .writedata
			audio_out_data_audio_s1_chipselect              => mm_interconnect_0_audio_out_data_audio_s1_chipselect,      --                                          .chipselect
			audio_out_pause_s1_address                      => mm_interconnect_0_audio_out_pause_s1_address,              --                        audio_out_pause_s1.address
			audio_out_pause_s1_write                        => mm_interconnect_0_audio_out_pause_s1_write,                --                                          .write
			audio_out_pause_s1_readdata                     => mm_interconnect_0_audio_out_pause_s1_readdata,             --                                          .readdata
			audio_out_pause_s1_writedata                    => mm_interconnect_0_audio_out_pause_s1_writedata,            --                                          .writedata
			audio_out_pause_s1_chipselect                   => mm_interconnect_0_audio_out_pause_s1_chipselect,           --                                          .chipselect
			audio_out_stop_s1_address                       => mm_interconnect_0_audio_out_stop_s1_address,               --                         audio_out_stop_s1.address
			audio_out_stop_s1_write                         => mm_interconnect_0_audio_out_stop_s1_write,                 --                                          .write
			audio_out_stop_s1_readdata                      => mm_interconnect_0_audio_out_stop_s1_readdata,              --                                          .readdata
			audio_out_stop_s1_writedata                     => mm_interconnect_0_audio_out_stop_s1_writedata,             --                                          .writedata
			audio_out_stop_s1_chipselect                    => mm_interconnect_0_audio_out_stop_s1_chipselect,            --                                          .chipselect
			audio_wrclk_s1_address                          => mm_interconnect_0_audio_wrclk_s1_address,                  --                            audio_wrclk_s1.address
			audio_wrclk_s1_write                            => mm_interconnect_0_audio_wrclk_s1_write,                    --                                          .write
			audio_wrclk_s1_readdata                         => mm_interconnect_0_audio_wrclk_s1_readdata,                 --                                          .readdata
			audio_wrclk_s1_writedata                        => mm_interconnect_0_audio_wrclk_s1_writedata,                --                                          .writedata
			audio_wrclk_s1_chipselect                       => mm_interconnect_0_audio_wrclk_s1_chipselect,               --                                          .chipselect
			audio_wrreq_s1_address                          => mm_interconnect_0_audio_wrreq_s1_address,                  --                            audio_wrreq_s1.address
			audio_wrreq_s1_write                            => mm_interconnect_0_audio_wrreq_s1_write,                    --                                          .write
			audio_wrreq_s1_readdata                         => mm_interconnect_0_audio_wrreq_s1_readdata,                 --                                          .readdata
			audio_wrreq_s1_writedata                        => mm_interconnect_0_audio_wrreq_s1_writedata,                --                                          .writedata
			audio_wrreq_s1_chipselect                       => mm_interconnect_0_audio_wrreq_s1_chipselect,               --                                          .chipselect
			audio_sel_s1_address                            => mm_interconnect_0_audio_sel_s1_address,                    --                              audio_sel_s1.address
			audio_sel_s1_write                              => mm_interconnect_0_audio_sel_s1_write,                      --                                          .write
			audio_sel_s1_readdata                           => mm_interconnect_0_audio_sel_s1_readdata,                   --                                          .readdata
			audio_sel_s1_writedata                          => mm_interconnect_0_audio_sel_s1_writedata,                  --                                          .writedata
			audio_sel_s1_chipselect                         => mm_interconnect_0_audio_sel_s1_chipselect,                 --                                          .chipselect
			cpu_jtag_debug_module_address                   => mm_interconnect_0_cpu_jtag_debug_module_address,           --                     cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write                     => mm_interconnect_0_cpu_jtag_debug_module_write,             --                                          .write
			cpu_jtag_debug_module_read                      => mm_interconnect_0_cpu_jtag_debug_module_read,              --                                          .read
			cpu_jtag_debug_module_readdata                  => mm_interconnect_0_cpu_jtag_debug_module_readdata,          --                                          .readdata
			cpu_jtag_debug_module_writedata                 => mm_interconnect_0_cpu_jtag_debug_module_writedata,         --                                          .writedata
			cpu_jtag_debug_module_byteenable                => mm_interconnect_0_cpu_jtag_debug_module_byteenable,        --                                          .byteenable
			cpu_jtag_debug_module_waitrequest               => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,       --                                          .waitrequest
			cpu_jtag_debug_module_debugaccess               => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,       --                                          .debugaccess
			dds_increment_s1_address                        => mm_interconnect_0_dds_increment_s1_address,                --                          dds_increment_s1.address
			dds_increment_s1_write                          => mm_interconnect_0_dds_increment_s1_write,                  --                                          .write
			dds_increment_s1_readdata                       => mm_interconnect_0_dds_increment_s1_readdata,               --                                          .readdata
			dds_increment_s1_writedata                      => mm_interconnect_0_dds_increment_s1_writedata,              --                                          .writedata
			dds_increment_s1_chipselect                     => mm_interconnect_0_dds_increment_s1_chipselect,             --                                          .chipselect
			div_freq_s1_address                             => mm_interconnect_0_div_freq_s1_address,                     --                               div_freq_s1.address
			div_freq_s1_write                               => mm_interconnect_0_div_freq_s1_write,                       --                                          .write
			div_freq_s1_readdata                            => mm_interconnect_0_div_freq_s1_readdata,                    --                                          .readdata
			div_freq_s1_writedata                           => mm_interconnect_0_div_freq_s1_writedata,                   --                                          .writedata
			div_freq_s1_chipselect                          => mm_interconnect_0_div_freq_s1_chipselect,                  --                                          .chipselect
			jtag_uart_avalon_jtag_slave_address             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --               jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                          .write
			jtag_uart_avalon_jtag_slave_read                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                          .read
			jtag_uart_avalon_jtag_slave_readdata            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                          .readdata
			jtag_uart_avalon_jtag_slave_writedata           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                          .writedata
			jtag_uart_avalon_jtag_slave_waitrequest         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                          .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                          .chipselect
			key_s1_address                                  => mm_interconnect_0_key_s1_address,                          --                                    key_s1.address
			key_s1_write                                    => mm_interconnect_0_key_s1_write,                            --                                          .write
			key_s1_readdata                                 => mm_interconnect_0_key_s1_readdata,                         --                                          .readdata
			key_s1_writedata                                => mm_interconnect_0_key_s1_writedata,                        --                                          .writedata
			key_s1_chipselect                               => mm_interconnect_0_key_s1_chipselect,                       --                                          .chipselect
			keyboard_keys_s1_address                        => mm_interconnect_0_keyboard_keys_s1_address,                --                          keyboard_keys_s1.address
			keyboard_keys_s1_readdata                       => mm_interconnect_0_keyboard_keys_s1_readdata,               --                                          .readdata
			lfsr_clk_interrupt_gen_s1_address               => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_address,       --                 lfsr_clk_interrupt_gen_s1.address
			lfsr_clk_interrupt_gen_s1_write                 => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write,         --                                          .write
			lfsr_clk_interrupt_gen_s1_readdata              => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_readdata,      --                                          .readdata
			lfsr_clk_interrupt_gen_s1_writedata             => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_writedata,     --                                          .writedata
			lfsr_clk_interrupt_gen_s1_chipselect            => mm_interconnect_0_lfsr_clk_interrupt_gen_s1_chipselect,    --                                          .chipselect
			lfsr_val_s1_address                             => mm_interconnect_0_lfsr_val_s1_address,                     --                               lfsr_val_s1.address
			lfsr_val_s1_readdata                            => mm_interconnect_0_lfsr_val_s1_readdata,                    --                                          .readdata
			modulation_selector_s1_address                  => mm_interconnect_0_modulation_selector_s1_address,          --                    modulation_selector_s1.address
			modulation_selector_s1_write                    => mm_interconnect_0_modulation_selector_s1_write,            --                                          .write
			modulation_selector_s1_readdata                 => mm_interconnect_0_modulation_selector_s1_readdata,         --                                          .readdata
			modulation_selector_s1_writedata                => mm_interconnect_0_modulation_selector_s1_writedata,        --                                          .writedata
			modulation_selector_s1_chipselect               => mm_interconnect_0_modulation_selector_s1_chipselect,       --                                          .chipselect
			mouse_pos_s1_address                            => mm_interconnect_0_mouse_pos_s1_address,                    --                              mouse_pos_s1.address
			mouse_pos_s1_readdata                           => mm_interconnect_0_mouse_pos_s1_readdata,                   --                                          .readdata
			sdram_s1_address                                => mm_interconnect_0_sdram_s1_address,                        --                                  sdram_s1.address
			sdram_s1_write                                  => mm_interconnect_0_sdram_s1_write,                          --                                          .write
			sdram_s1_read                                   => mm_interconnect_0_sdram_s1_read,                           --                                          .read
			sdram_s1_readdata                               => mm_interconnect_0_sdram_s1_readdata,                       --                                          .readdata
			sdram_s1_writedata                              => mm_interconnect_0_sdram_s1_writedata,                      --                                          .writedata
			sdram_s1_byteenable                             => mm_interconnect_0_sdram_s1_byteenable,                     --                                          .byteenable
			sdram_s1_readdatavalid                          => mm_interconnect_0_sdram_s1_readdatavalid,                  --                                          .readdatavalid
			sdram_s1_waitrequest                            => mm_interconnect_0_sdram_s1_waitrequest,                    --                                          .waitrequest
			sdram_s1_chipselect                             => mm_interconnect_0_sdram_s1_chipselect,                     --                                          .chipselect
			signal_selector_s1_address                      => mm_interconnect_0_signal_selector_s1_address,              --                        signal_selector_s1.address
			signal_selector_s1_write                        => mm_interconnect_0_signal_selector_s1_write,                --                                          .write
			signal_selector_s1_readdata                     => mm_interconnect_0_signal_selector_s1_readdata,             --                                          .readdata
			signal_selector_s1_writedata                    => mm_interconnect_0_signal_selector_s1_writedata,            --                                          .writedata
			signal_selector_s1_chipselect                   => mm_interconnect_0_signal_selector_s1_chipselect,           --                                          .chipselect
			sysid_qsys_control_slave_address                => mm_interconnect_0_sysid_qsys_control_slave_address,        --                  sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata               => mm_interconnect_0_sysid_qsys_control_slave_readdata,       --                                          .readdata
			timer_s1_address                                => mm_interconnect_0_timer_s1_address,                        --                                  timer_s1.address
			timer_s1_write                                  => mm_interconnect_0_timer_s1_write,                          --                                          .write
			timer_s1_readdata                               => mm_interconnect_0_timer_s1_readdata,                       --                                          .readdata
			timer_s1_writedata                              => mm_interconnect_0_timer_s1_writedata,                      --                                          .writedata
			timer_s1_chipselect                             => mm_interconnect_0_timer_s1_chipselect,                     --                                          .chipselect
			vga_to_nios_2_datamaster_address                => mm_interconnect_0_vga_to_nios_2_datamaster_address,        --                  vga_to_nios_2_datamaster.address
			vga_to_nios_2_datamaster_write                  => mm_interconnect_0_vga_to_nios_2_datamaster_write,          --                                          .write
			vga_to_nios_2_datamaster_read                   => mm_interconnect_0_vga_to_nios_2_datamaster_read,           --                                          .read
			vga_to_nios_2_datamaster_readdata               => mm_interconnect_0_vga_to_nios_2_datamaster_readdata,       --                                          .readdata
			vga_to_nios_2_datamaster_writedata              => mm_interconnect_0_vga_to_nios_2_datamaster_writedata       --                                          .writedata
		);

	irq_mapper : component DE1_SoC_QSYS_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			sender_irq    => cpu_d_irq_irq                       --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk0_clk,                    --       receiver_clk.clk
			sender_clk     => clk_clk,                            --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_002_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	rst_controller : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => pll_outclk0_clk,                --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component de1_soc_qsys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,      -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_outclk2_clk,                    --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => vga_vga_clk_clk_internal,           --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_audio_data_fregen_s1_write_ports_inv <= not mm_interconnect_0_audio_data_fregen_s1_write;

	mm_interconnect_0_audio_out_data_audio_s1_write_ports_inv <= not mm_interconnect_0_audio_out_data_audio_s1_write;

	mm_interconnect_0_audio_out_pause_s1_write_ports_inv <= not mm_interconnect_0_audio_out_pause_s1_write;

	mm_interconnect_0_audio_out_stop_s1_write_ports_inv <= not mm_interconnect_0_audio_out_stop_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_signal_selector_s1_write_ports_inv <= not mm_interconnect_0_signal_selector_s1_write;

	mm_interconnect_0_modulation_selector_s1_write_ports_inv <= not mm_interconnect_0_modulation_selector_s1_write;

	mm_interconnect_0_div_freq_s1_write_ports_inv <= not mm_interconnect_0_div_freq_s1_write;

	mm_interconnect_0_audio_sel_s1_write_ports_inv <= not mm_interconnect_0_audio_sel_s1_write;

	mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write_ports_inv <= not mm_interconnect_0_lfsr_clk_interrupt_gen_s1_write;

	mm_interconnect_0_dds_increment_s1_write_ports_inv <= not mm_interconnect_0_dds_increment_s1_write;

	mm_interconnect_0_audio_wrclk_s1_write_ports_inv <= not mm_interconnect_0_audio_wrclk_s1_write;

	mm_interconnect_0_audio_wrreq_s1_write_ports_inv <= not mm_interconnect_0_audio_wrreq_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	clk_25_out_clk <= pll_outclk2_clk;

	vga_vga_clk_clk <= vga_vga_clk_clk_internal;

end architecture rtl; -- of DE1_SoC_QSYS
