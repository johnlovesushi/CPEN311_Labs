module DDS ( input clk,
				 input  [31:0] in,
				 output [11:0] out);
	
endmodule
