-- DE1_SoC_QSYS_vga.vhd

-- Generated using ACDS version 14.1 186 at 2017.11.28.14:39:07

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE1_SoC_QSYS_vga is
	port (
		alt_vip_itc_0_clocked_video_vid_clk       : in  std_logic                     := '0';             --    alt_vip_itc_0_clocked_video.vid_clk
		alt_vip_itc_0_clocked_video_vid_data      : out std_logic_vector(23 downto 0);                    --                               .vid_data
		alt_vip_itc_0_clocked_video_underflow     : out std_logic;                                        --                               .underflow
		alt_vip_itc_0_clocked_video_vid_datavalid : out std_logic;                                        --                               .vid_datavalid
		alt_vip_itc_0_clocked_video_vid_v_sync    : out std_logic;                                        --                               .vid_v_sync
		alt_vip_itc_0_clocked_video_vid_h_sync    : out std_logic;                                        --                               .vid_h_sync
		alt_vip_itc_0_clocked_video_vid_f         : out std_logic;                                        --                               .vid_f
		alt_vip_itc_0_clocked_video_vid_h         : out std_logic;                                        --                               .vid_h
		alt_vip_itc_0_clocked_video_vid_v         : out std_logic;                                        --                               .vid_v
		alt_vip_vfr_0_interrupt_sender_irq        : out std_logic;                                        -- alt_vip_vfr_0_interrupt_sender.irq
		clk_50m_clk                               : in  std_logic                     := '0';             --                        clk_50m.clk
		clk_50m_reset_reset_n                     : in  std_logic                     := '0';             --                  clk_50m_reset.reset_n
		nios_clk_clk                              : in  std_logic                     := '0';             --                       nios_clk.clk
		nios_clk_reset_reset_n                    : in  std_logic                     := '0';             --                 nios_clk_reset.reset_n
		to_nios_2_datamaster_address              : in  std_logic_vector(4 downto 0)  := (others => '0'); --           to_nios_2_datamaster.address
		to_nios_2_datamaster_write                : in  std_logic                     := '0';             --                               .write
		to_nios_2_datamaster_writedata            : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		to_nios_2_datamaster_read                 : in  std_logic                     := '0';             --                               .read
		to_nios_2_datamaster_readdata             : out std_logic_vector(31 downto 0);                    --                               .readdata
		to_sdram_address                          : out std_logic_vector(31 downto 0);                    --                       to_sdram.address
		to_sdram_burstcount                       : out std_logic_vector(5 downto 0);                     --                               .burstcount
		to_sdram_readdata                         : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .readdata
		to_sdram_read                             : out std_logic;                                        --                               .read
		to_sdram_readdatavalid                    : in  std_logic                     := '0';             --                               .readdatavalid
		to_sdram_waitrequest                      : in  std_logic                     := '0';             --                               .waitrequest
		vga_clk_clk                               : out std_logic                                         --                        vga_clk.clk
	);
end entity DE1_SoC_QSYS_vga;

architecture rtl of DE1_SoC_QSYS_vga is
	component alt_vipitc131_IS2Vid is
		generic (
			NUMBER_OF_COLOUR_PLANES       : integer := 3;
			COLOUR_PLANES_ARE_IN_PARALLEL : integer := 1;
			BPS                           : integer := 8;
			INTERLACED                    : integer := 0;
			H_ACTIVE_PIXELS               : integer := 1920;
			V_ACTIVE_LINES                : integer := 1200;
			ACCEPT_COLOURS_IN_SEQ         : integer := 0;
			FIFO_DEPTH                    : integer := 1920;
			CLOCKS_ARE_SAME               : integer := 0;
			USE_CONTROL                   : integer := 0;
			NO_OF_MODES                   : integer := 1;
			THRESHOLD                     : integer := 1919;
			STD_WIDTH                     : integer := 1;
			GENERATE_SYNC                 : integer := 0;
			USE_EMBEDDED_SYNCS            : integer := 0;
			AP_LINE                       : integer := 0;
			V_BLANK                       : integer := 0;
			H_BLANK                       : integer := 0;
			H_SYNC_LENGTH                 : integer := 44;
			H_FRONT_PORCH                 : integer := 88;
			H_BACK_PORCH                  : integer := 148;
			V_SYNC_LENGTH                 : integer := 5;
			V_FRONT_PORCH                 : integer := 4;
			V_BACK_PORCH                  : integer := 36;
			F_RISING_EDGE                 : integer := 0;
			F_FALLING_EDGE                : integer := 0;
			FIELD0_V_RISING_EDGE          : integer := 0;
			FIELD0_V_BLANK                : integer := 0;
			FIELD0_V_SYNC_LENGTH          : integer := 0;
			FIELD0_V_FRONT_PORCH          : integer := 0;
			FIELD0_V_BACK_PORCH           : integer := 0;
			ANC_LINE                      : integer := 0;
			FIELD0_ANC_LINE               : integer := 0
		);
		port (
			is_clk        : in  std_logic                     := 'X';             -- clk
			rst           : in  std_logic                     := 'X';             -- reset
			is_data       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			is_valid      : in  std_logic                     := 'X';             -- valid
			is_ready      : out std_logic;                                        -- ready
			is_sop        : in  std_logic                     := 'X';             -- startofpacket
			is_eop        : in  std_logic                     := 'X';             -- endofpacket
			vid_clk       : in  std_logic                     := 'X';             -- export
			vid_data      : out std_logic_vector(23 downto 0);                    -- export
			underflow     : out std_logic;                                        -- export
			vid_datavalid : out std_logic;                                        -- export
			vid_v_sync    : out std_logic;                                        -- export
			vid_h_sync    : out std_logic;                                        -- export
			vid_f         : out std_logic;                                        -- export
			vid_h         : out std_logic;                                        -- export
			vid_v         : out std_logic                                         -- export
		);
	end component alt_vipitc131_IS2Vid;

	component alt_vipvfr131_vfr is
		generic (
			BITS_PER_PIXEL_PER_COLOR_PLANE : integer := 8;
			NUMBER_OF_CHANNELS_IN_PARALLEL : integer := 3;
			NUMBER_OF_CHANNELS_IN_SEQUENCE : integer := 1;
			MAX_IMAGE_WIDTH                : integer := 640;
			MAX_IMAGE_HEIGHT               : integer := 480;
			MEM_PORT_WIDTH                 : integer := 256;
			RMASTER_FIFO_DEPTH             : integer := 64;
			RMASTER_BURST_TARGET           : integer := 32;
			CLOCKS_ARE_SEPARATE            : integer := 1
		);
		port (
			clock                : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_clock         : in  std_logic                     := 'X';             -- clk
			master_reset         : in  std_logic                     := 'X';             -- reset
			slave_address        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			slave_irq            : out std_logic;                                        -- irq
			dout_data            : out std_logic_vector(23 downto 0);                    -- data
			dout_valid           : out std_logic;                                        -- valid
			dout_ready           : in  std_logic                     := 'X';             -- ready
			dout_startofpacket   : out std_logic;                                        -- startofpacket
			dout_endofpacket     : out std_logic;                                        -- endofpacket
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_burstcount    : out std_logic_vector(5 downto 0);                     -- burstcount
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X'              -- waitrequest
		);
	end component alt_vipvfr131_vfr;

	component DE1_SoC_QSYS_vga_vga_clk is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DE1_SoC_QSYS_vga_vga_clk;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal alt_vip_vfr_0_avalon_streaming_source_valid         : std_logic;                     -- alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	signal alt_vip_vfr_0_avalon_streaming_source_data          : std_logic_vector(23 downto 0); -- alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	signal alt_vip_vfr_0_avalon_streaming_source_ready         : std_logic;                     -- alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	signal alt_vip_vfr_0_avalon_streaming_source_startofpacket : std_logic;                     -- alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	signal alt_vip_vfr_0_avalon_streaming_source_endofpacket   : std_logic;                     -- alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	signal rst_controller_reset_out_reset                      : std_logic;                     -- rst_controller:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_0:master_reset, alt_vip_vfr_0:reset]
	signal clk_50m_reset_reset_n_ports_inv                     : std_logic;                     -- clk_50m_reset_reset_n:inv -> vga_clk:rst
	signal nios_clk_reset_reset_n_ports_inv                    : std_logic;                     -- nios_clk_reset_reset_n:inv -> rst_controller:reset_in0

begin

	alt_vip_itc_0 : component alt_vipitc131_IS2Vid
		generic map (
			NUMBER_OF_COLOUR_PLANES       => 3,
			COLOUR_PLANES_ARE_IN_PARALLEL => 1,
			BPS                           => 8,
			INTERLACED                    => 0,
			H_ACTIVE_PIXELS               => 800,
			V_ACTIVE_LINES                => 600,
			ACCEPT_COLOURS_IN_SEQ         => 0,
			FIFO_DEPTH                    => 512,
			CLOCKS_ARE_SAME               => 0,
			USE_CONTROL                   => 0,
			NO_OF_MODES                   => 1,
			THRESHOLD                     => 450,
			STD_WIDTH                     => 1,
			GENERATE_SYNC                 => 0,
			USE_EMBEDDED_SYNCS            => 0,
			AP_LINE                       => 0,
			V_BLANK                       => 0,
			H_BLANK                       => 0,
			H_SYNC_LENGTH                 => 128,
			H_FRONT_PORCH                 => 40,
			H_BACK_PORCH                  => 88,
			V_SYNC_LENGTH                 => 4,
			V_FRONT_PORCH                 => 1,
			V_BACK_PORCH                  => 23,
			F_RISING_EDGE                 => 0,
			F_FALLING_EDGE                => 0,
			FIELD0_V_RISING_EDGE          => 0,
			FIELD0_V_BLANK                => 0,
			FIELD0_V_SYNC_LENGTH          => 0,
			FIELD0_V_FRONT_PORCH          => 0,
			FIELD0_V_BACK_PORCH           => 0,
			ANC_LINE                      => 0,
			FIELD0_ANC_LINE               => 0
		)
		port map (
			is_clk        => nios_clk_clk,                                        --       is_clk_rst.clk
			rst           => rst_controller_reset_out_reset,                      -- is_clk_rst_reset.reset
			is_data       => alt_vip_vfr_0_avalon_streaming_source_data,          --              din.data
			is_valid      => alt_vip_vfr_0_avalon_streaming_source_valid,         --                 .valid
			is_ready      => alt_vip_vfr_0_avalon_streaming_source_ready,         --                 .ready
			is_sop        => alt_vip_vfr_0_avalon_streaming_source_startofpacket, --                 .startofpacket
			is_eop        => alt_vip_vfr_0_avalon_streaming_source_endofpacket,   --                 .endofpacket
			vid_clk       => alt_vip_itc_0_clocked_video_vid_clk,                 --    clocked_video.export
			vid_data      => alt_vip_itc_0_clocked_video_vid_data,                --                 .export
			underflow     => alt_vip_itc_0_clocked_video_underflow,               --                 .export
			vid_datavalid => alt_vip_itc_0_clocked_video_vid_datavalid,           --                 .export
			vid_v_sync    => alt_vip_itc_0_clocked_video_vid_v_sync,              --                 .export
			vid_h_sync    => alt_vip_itc_0_clocked_video_vid_h_sync,              --                 .export
			vid_f         => alt_vip_itc_0_clocked_video_vid_f,                   --                 .export
			vid_h         => alt_vip_itc_0_clocked_video_vid_h,                   --                 .export
			vid_v         => alt_vip_itc_0_clocked_video_vid_v                    --                 .export
		);

	alt_vip_vfr_0 : component alt_vipvfr131_vfr
		generic map (
			BITS_PER_PIXEL_PER_COLOR_PLANE => 8,
			NUMBER_OF_CHANNELS_IN_PARALLEL => 3,
			NUMBER_OF_CHANNELS_IN_SEQUENCE => 1,
			MAX_IMAGE_WIDTH                => 800,
			MAX_IMAGE_HEIGHT               => 600,
			MEM_PORT_WIDTH                 => 32,
			RMASTER_FIFO_DEPTH             => 64,
			RMASTER_BURST_TARGET           => 32,
			CLOCKS_ARE_SEPARATE            => 1
		)
		port map (
			clock                => nios_clk_clk,                                        --             clock_reset.clk
			reset                => rst_controller_reset_out_reset,                      --       clock_reset_reset.reset
			master_clock         => nios_clk_clk,                                        --            clock_master.clk
			master_reset         => rst_controller_reset_out_reset,                      --      clock_master_reset.reset
			slave_address        => to_nios_2_datamaster_address,                        --            avalon_slave.address
			slave_write          => to_nios_2_datamaster_write,                          --                        .write
			slave_writedata      => to_nios_2_datamaster_writedata,                      --                        .writedata
			slave_read           => to_nios_2_datamaster_read,                           --                        .read
			slave_readdata       => to_nios_2_datamaster_readdata,                       --                        .readdata
			slave_irq            => alt_vip_vfr_0_interrupt_sender_irq,                  --        interrupt_sender.irq
			dout_data            => alt_vip_vfr_0_avalon_streaming_source_data,          -- avalon_streaming_source.data
			dout_valid           => alt_vip_vfr_0_avalon_streaming_source_valid,         --                        .valid
			dout_ready           => alt_vip_vfr_0_avalon_streaming_source_ready,         --                        .ready
			dout_startofpacket   => alt_vip_vfr_0_avalon_streaming_source_startofpacket, --                        .startofpacket
			dout_endofpacket     => alt_vip_vfr_0_avalon_streaming_source_endofpacket,   --                        .endofpacket
			master_address       => to_sdram_address,                                    --           avalon_master.address
			master_burstcount    => to_sdram_burstcount,                                 --                        .burstcount
			master_readdata      => to_sdram_readdata,                                   --                        .readdata
			master_read          => to_sdram_read,                                       --                        .read
			master_readdatavalid => to_sdram_readdatavalid,                              --                        .readdatavalid
			master_waitrequest   => to_sdram_waitrequest                                 --                        .waitrequest
		);

	vga_clk : component DE1_SoC_QSYS_vga_vga_clk
		port map (
			refclk   => clk_50m_clk,                     --  refclk.clk
			rst      => clk_50m_reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => vga_clk_clk,                     -- outclk0.clk
			locked   => open                             -- (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios_clk_reset_reset_n_ports_inv, -- reset_in0.reset
			clk            => nios_clk_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                             -- (terminated)
			reset_req_in0  => '0',                              -- (terminated)
			reset_in1      => '0',                              -- (terminated)
			reset_req_in1  => '0',                              -- (terminated)
			reset_in2      => '0',                              -- (terminated)
			reset_req_in2  => '0',                              -- (terminated)
			reset_in3      => '0',                              -- (terminated)
			reset_req_in3  => '0',                              -- (terminated)
			reset_in4      => '0',                              -- (terminated)
			reset_req_in4  => '0',                              -- (terminated)
			reset_in5      => '0',                              -- (terminated)
			reset_req_in5  => '0',                              -- (terminated)
			reset_in6      => '0',                              -- (terminated)
			reset_req_in6  => '0',                              -- (terminated)
			reset_in7      => '0',                              -- (terminated)
			reset_req_in7  => '0',                              -- (terminated)
			reset_in8      => '0',                              -- (terminated)
			reset_req_in8  => '0',                              -- (terminated)
			reset_in9      => '0',                              -- (terminated)
			reset_req_in9  => '0',                              -- (terminated)
			reset_in10     => '0',                              -- (terminated)
			reset_req_in10 => '0',                              -- (terminated)
			reset_in11     => '0',                              -- (terminated)
			reset_req_in11 => '0',                              -- (terminated)
			reset_in12     => '0',                              -- (terminated)
			reset_req_in12 => '0',                              -- (terminated)
			reset_in13     => '0',                              -- (terminated)
			reset_req_in13 => '0',                              -- (terminated)
			reset_in14     => '0',                              -- (terminated)
			reset_req_in14 => '0',                              -- (terminated)
			reset_in15     => '0',                              -- (terminated)
			reset_req_in15 => '0'                               -- (terminated)
		);

	clk_50m_reset_reset_n_ports_inv <= not clk_50m_reset_reset_n;

	nios_clk_reset_reset_n_ports_inv <= not nios_clk_reset_reset_n;

end architecture rtl; -- of DE1_SoC_QSYS_vga
